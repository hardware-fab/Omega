//----------------------------------------------------------------------------
//  This file is a part of the VESPA SoC Prototyping Framework
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the Apache 2.0 License.
//
// File:    bram36.vhd
// Authors: Gabriele Montanaro
//          Andrea Galimberti
//          Davide Zoni
// Company: Politecnico di Milano
// Mail:    name.surname@polimi.it
//
// ----------------------------------------------------------------------------

module bram36 #(
    parameter READ_WIDTH            = 36,
    parameter WRITE_WIDTH           = 36,
    parameter ADDR_WIDTH            = 10,
    parameter WE_WIDTH              = 4
    )
    (
    input                        clk,
    input                        reset,
    input  [ADDR_WIDTH-1:0]      addr_i,
    input                        valid_i,
    output [READ_WIDTH-1:0]      data_o
    );
    wire [WRITE_WIDTH-1:0] data_i ;
    wire [WE_WIDTH-1:0]    we ;
    wire                   regce;
    assign  we      = { WE_WIDTH{1'b0}    };
    assign  data_i  = { WRITE_WIDTH{1'b0} };
    assign  regce   = 1'b0;
    BRAM_SINGLE_MACRO #(
        .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
        .DEVICE("7SERIES"), // Target Device: "7SERIES" 
        .DO_REG(0), // Optional output register (0 or 1)
        .INIT(36'b000000000000000000000000000000000000), // Initial values on output port
        .INIT_FILE ("NONE"),
        .WRITE_WIDTH(WRITE_WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(READ_WIDTH),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .SRVAL(36'b000000000000000000000000000000000000), // Set/Reset value for port output
        .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        .INIT_00(256'h00080440000704400006044000060480000604e000060580000605c000060780),
.INIT_01(256'h010804a001060480010704a0000604a0000604a0000b0440000604c000090440),
.INIT_02(256'h0206046001060460010604600106046001060460010904a0010904a0010804a0),
.INIT_03(256'h0206046002060460020604600206046002060460020604600206046002060460),
.INIT_04(256'h0306046003060460030604600306046003060460030604600306046002060460),
.INIT_05(256'h0406046004060460040604600406046004060460030604600306046003060460),
.INIT_06(256'h0506046005060460050604600406046004060460040604600406046004060460),
.INIT_07(256'h0606046005060460050604600506046005060460050604600506046005060460),
.INIT_08(256'h0606046006060460060604600606046006060460060604600606046006060460),
.INIT_09(256'h0706046007060460070604600706046007060460070604600706046006060460),
.INIT_0A(256'h0806046008060460080604600806046008060460070604600706046007060460),
.INIT_0B(256'h0906046009060460090604600806046008060460080604600806046008060460),
.INIT_0C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_0D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_0E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_0F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_10(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_11(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_12(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_13(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_14(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_15(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_16(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_17(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_18(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_19(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_1F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_20(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_21(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_22(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_23(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_24(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_25(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_26(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_27(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_28(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_29(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_2F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_30(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_31(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_32(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_33(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_34(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_35(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_36(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_37(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_38(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_39(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_3F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_40(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_41(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_42(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_43(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_44(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_45(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_46(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_47(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_48(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_49(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_4F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_50(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_51(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_52(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_53(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_54(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_55(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_56(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_57(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_58(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_59(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_5F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_60(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_61(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_62(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_63(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_64(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_65(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_66(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_67(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_68(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_69(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_6F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_70(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_71(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_72(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_73(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_74(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_75(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_76(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_77(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_78(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_79(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7A(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7B(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7C(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7D(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7E(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INIT_7F(256'h0906046009060460090604600906046009060460090604600906046009060460),
.INITP_00(256'h0444440000044444000004444400000444440000044446020006454511111011),
.INITP_01(256'h4444444444444444444444444444440000044444000004444400000444440000),
.INITP_02(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_03(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_04(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_05(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_06(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_07(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_08(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_09(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0A(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0B(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0C(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0D(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0E(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0F(256'h4444444444444444444444444444444444444444444444444444444444444444)) 
        BRAM_SINGLE_MACRO_inst (
            .DO(data_o),   // Output data, width defined by READ_WIDTH parameter
            .ADDR(addr_i), // Input address, width defined by read/write port depth look at the table below
            .CLK(clk),     // 1-bit input clock
            .DI(data_i),   // Input data port, width defined by WRITE_WIDTH parameter
            .EN(valid_i),  // 1-bit input RAM enable
            .REGCE(regce), // 1-bit input output register enable
            .RST(reset),   // 1-bit input reset
            .WE(we)        // Input write enable, width defined by write port depth look at tabel below
        );
        /////////////////////////////////////////////////////////////////////
        //  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            //
        // WRITE_WIDTH |           | WRITE Depth |            |  WE Width  //
        // ============|===========|=============|============|============//
        //    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   //
        //    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   //
        //    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   //
        //    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   //
        //    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   //
        //     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   //
        //     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   //
        //     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   //
        //     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   //
        //       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   //
        //       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   //
        //       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   //
        //       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   //
        /////////////////////////////////////////////////////////////////////
        
 endmodule
