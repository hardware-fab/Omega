//----------------------------------------------------------------------------
//  This file is a part of the VESPA SoC Prototyping Framework
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the Apache 2.0 License.
//
// File:    bram36_old.vhd
// Authors: Gabriele Montanaro
//          Andrea Galimberti
//          Davide Zoni
// Company: Politecnico di Milano
// Mail:    name.surname@polimi.it
//
// ----------------------------------------------------------------------------

module bram36 #(
    parameter READ_WIDTH            = 36,
    parameter WRITE_WIDTH           = 36,
    parameter ADDR_WIDTH            = 10,
    parameter WE_WIDTH              = 4
    )
    (
    input                        clk,
    input                        reset,
    input  [ADDR_WIDTH-1:0]      addr_i,
    input                        valid_i,
    output [READ_WIDTH-1:0]      data_o
    );
    wire [WRITE_WIDTH-1:0] data_i ;
    wire [WE_WIDTH-1:0]    we ;
    wire                   regce;
    assign  we      = { WE_WIDTH{1'b0}    };
    assign  data_i  = { WRITE_WIDTH{1'b0} };
    assign  regce   = 1'b0;
    BRAM_SINGLE_MACRO #(
        .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
        .DEVICE("7SERIES"), // Target Device: "7SERIES" 
        .DO_REG(0), // Optional output register (0 or 1)
        .INIT(36'b000000000000000000000000000000000000), // Initial values on output port
        .INIT_FILE ("NONE"),
        .WRITE_WIDTH(WRITE_WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(READ_WIDTH),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .SRVAL(36'b000000000000000000000000000000000000), // Set/Reset value for port output
        .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        .INIT_00(256'h000f08d6000604b200090416000604c0000604ea00060440000604e0000605c0),
.INIT_01(256'h000904da000604a0000b0416000e08b2000e08ba000704b2000b0440000d08b2),
.INIT_02(256'h0007049e000804b2000b04ee000804be000604a0000804b2000b040a000f08b2),
.INIT_03(256'h010804c0010e088a01060472010c087e010c087e010b04ee010804a6000704a0),
.INIT_04(256'h010b0400010a04d60106046e0107049201070492010f089e010c04fe010c04fe),
.INIT_05(256'h020f08960206046a0206046a010e08a0010a04d20107048e010f089a010904b2),
.INIT_06(256'h04060466040904be030a04ca030c0872020c04ee0206047e0207048a020a04ce),
.INIT_07(256'h08060480080f088e070c086e070904ba060a04c6060904a605070486050b04de),
.INIT_08(256'h106b04d20c6c086a0b0f088a0b0f088a0a0604760a0904b6090b04d609060480),
.INIT_09(256'h306c08662c6904ae286f0886246b04ce206604721c68049218680492146904b2),
.INIT_0A(256'h506b04c64c6a04be4866046e446f08a0406b04de3c6b04ca3868048e346c0866),
.INIT_0B(256'h7067047e6c66046a686b04d6646a04ba606904a65c6d0876586c0880546b04da),
.INIT_0C(256'h8306046683060466830d0872830d0872806d08727c6a04b6786904c074680486),
.INIT_0D(256'h830a04ae830b04ca830d086e830d086e830d086e830604668306046683060466),
.INIT_0E(256'h8308048e830e087e830a04aa830a04be830c04da830604808307047683080492),
.INIT_0F(256'h830e087a8309049e8309049e830a04a68307047283070472830b04e0830c04d6),
.INIT_10(256'h830804868309049a8307046e830c04ce830a04c0830a04b6830a04b68308048a),
.INIT_11(256'h8307046a83090496830904968307047e830d0880830c04ca830e0876830a04b2),
.INIT_12(256'h8307047a8307047a8307047a830b04be830b04be830e0872830804a0830804a0),
.INIT_13(256'h830704768309048e830a04a6830e086e830b04ba830b04ba8307046683070466),
.INIT_14(256'h830e086a8309048a83070480830704808309049e8306045e830b04b683070476),
.INIT_15(256'h8306045a8306045a830f087a830f087a8309049a8307047283070472830b04b2),
.INIT_16(256'h830f0876830b04aa8307046e8307046e83090496830e0866830e08668306045a),
.INIT_17(256'h8307046a830b04a6830e08808309049283090492830b04ba8308047e830904a0),
.INIT_18(256'h830a049e830b04c0830b04c08309048e8308047a830f0872830b04b6830b04b6),
.INIT_19(256'h830b04ae83080476830c085a830f086e8306045283060452830b04b2830b04b2),
.INIT_1A(256'h830b04aa830704808307048083070480830c04be830c04be830c04be830a049a),
.INIT_1B(256'h830b04a6830b04a68306045e8306045e830c0856830c08568306044e830f086a),
.INIT_1C(256'h830b04c08308047e8308046e8308046e830f0866830a0492830c04b6830904a0),
.INIT_1D(256'h830f0880830f0880830a049e830a049e830a048e8306045a830c08528306044a),
.INIT_1E(256'h83060446830a049a830a049a830a048a830a048a8308047a8308047a8308046a),
.INIT_1F(256'h830a0496830a0486830804768308046683080466830d085e83060456830c084e),
.INIT_20(256'h83060460830604608306046083060460830c04a6830c04a6830c04a6830c04a6),
.INIT_21(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_22(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_23(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_24(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_25(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_26(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_27(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_28(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_29(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_2F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_30(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_31(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_32(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_33(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_34(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_35(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_36(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_37(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_38(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_39(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_3F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_40(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_41(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_42(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_43(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_44(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_45(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_46(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_47(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_48(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_49(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_4F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_50(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_51(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_52(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_53(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_54(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_55(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_56(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_57(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_58(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_59(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_5F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_60(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_61(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_62(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_63(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_64(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_65(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_66(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_67(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_68(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_69(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_6F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_70(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_71(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_72(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_73(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_74(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_75(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_76(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_77(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_78(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_79(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7A(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7B(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7C(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7D(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7E(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INIT_7F(256'h8306046083060460830604608306046083060460830604608306046083060460),
.INITP_00(256'h4262606042624222200666647646620022022224664664764012201222302111),
.INITP_01(256'h6444446466464646466666666666202002202222002220022220200202626240),
.INITP_02(256'h6466664464666664446666646444644664664444666446664446646664444666),
.INITP_03(256'h6464466646644664666646646644644666666646666644446466446644464666),
.INITP_04(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_05(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_06(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_07(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_08(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_09(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0A(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0B(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0C(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0D(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0E(256'h4444444444444444444444444444444444444444444444444444444444444444),
.INITP_0F(256'h4444444444444444444444444444444444444444444444444444444444444444)) 
        BRAM_SINGLE_MACRO_inst (
            .DO(data_o),   // Output data, width defined by READ_WIDTH parameter
            .ADDR(addr_i), // Input address, width defined by read/write port depth look at the table below
            .CLK(clk),     // 1-bit input clock
            .DI(data_i),   // Input data port, width defined by WRITE_WIDTH parameter
            .EN(valid_i),  // 1-bit input RAM enable
            .REGCE(regce), // 1-bit input output register enable
            .RST(reset),   // 1-bit input reset
            .WE(we)        // Input write enable, width defined by write port depth look at tabel below
        );
        /////////////////////////////////////////////////////////////////////
        //  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            //
        // WRITE_WIDTH |           | WRITE Depth |            |  WE Width  //
        // ============|===========|=============|============|============//
        //    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   //
        //    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   //
        //    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   //
        //    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   //
        //    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   //
        //     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   //
        //     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   //
        //     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   //
        //     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   //
        //       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   //
        //       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   //
        //       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   //
        //       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   //
        /////////////////////////////////////////////////////////////////////
        
 endmodule
