-- Copyright (c) 2011-2023 Columbia University, System Level Design Group
-- SPDX-License-Identifier: Apache-2.0

------------------------------------------------------------------------------
--  ESP - xilinx - u55c
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


use work.grlib_config.all;
use work.amba.all;
use work.stdlib.all;
use work.devices.all;
use work.gencomp.all;
use work.leon3.all;
use work.uart.all;
use work.misc.all;
use work.net.all;
use work.svga_pkg.all;
library unisim;
-- pragma translate_off
use work.sim.all;
-- pragma translate_on
use unisim.VCOMPONENTS.all;
use work.monitor_pkg.all;
use work.sldacc.all;
use work.tile.all;
use work.nocpackage.all;
use work.cachepackage.all;
use work.coretypes.all;
use work.config.all;
use work.esp_global.all;
use work.socmap.all;
use work.tiles_pkg.all;

use work.esp_csr_pkg.all; --GM change: I need this library for freq data info
use work.hbm_pkg.all;


entity top is
  generic (
    SIMULATION          : boolean := false
  );
  port (
    clk_board_p            : in    std_ulogic;  -- 100 MHz clock
    clk_board_n            : in    std_ulogic;  -- 100 MHz clock
    --clk_hbm_p              : in    std_ulogic;  -- 100 MHz HBM reference clock 
    --clk_hbm_n              : in    std_ulogic;  -- 100 MHz HBM reference clock               
    cpu_reset_fpga         : in    std_ulogic;
    uart0_rxd              : in    std_ulogic;
    uart0_txd              : out   std_ulogic;
    dram_stat_catrip       : out   std_ulogic
    );
end;


architecture rtl of top is

--GM change: I add the declaration of the DFS module
component clockManager
  generic(
    PLL_FREQ                                 :    integer := 1;
    RANDOM_FREQ                              :    integer := 0
    --N_CLOCK_OUT                              :    integer := 1
  );
  port (
    rst_in                                   :     in std_logic;
    clk_in                                   :     in std_logic;
    mmcm_clk_o                               :     out std_ulogic;--_vector(N_CLOCK_OUT-1 downto 0);
    mmcm_locked_o                            :     out std_logic;
    freq_data_in                             :     in std_logic_vector(8-1 downto 0);
    freq_valid_in                            :     in std_logic
    );
end component;

function set_ddr_index (
  constant n : integer range 0 to 3)
  return integer is
begin
  if n > (MEM_ID_RANGE_MSB) then
    return MEM_ID_RANGE_MSB;
  else
    return n;
  end if;
end set_ddr_index;

constant this_ddr_index : attribute_vector(0 to 3) := (
  0 => set_ddr_index(0),
  1 => set_ddr_index(1),
  2 => set_ddr_index(2),
  3 => set_ddr_index(3)
  );

--Duration of the external reset pulse
constant EXT_RST_DURATION : integer := 100;

constant BAUDRATE         : positive := 38400;
constant BOARD_CLOCK_FREQ : positive := 100000000;
-------------------------------------------------------------------------------
-- Signals --------------------------------------------------------------------
-------------------------------------------------------------------------------

-- Clock and reset
signal clk_board              : std_ulogic;             --Clock generated by the u55c board. Freq: 100MHz
signal rst_board              : std_ulogic;             --Reset generated by the u55c board.
--signal clk_hbm                : std_ulogic;

signal sync_rst0, sync_rst1   : std_ulogic;             --Signals for the 2-stage flip-flop synchronizer for the input reset

signal clk_sys                : std_ulogic;             --Main system clock sent to the tiles
signal lock_sys               : std_ulogic;             --Lock signal of the main system clock

signal rstn_board             : std_ulogic;             --Negated profpga reset, synchronized with system clock
signal rstn_sys               : std_ulogic;             --Active low main system reset
signal rstn_init              : std_ulogic;             --Active low reset for clocking resources (synchronized with system clock)

signal cgi                    : clkgen_in_type;         --Clock generator input signal for the system clock
signal cgo                    : clkgen_out_type;        --Clock generator output signal for the system clock

signal lock_tiles             : std_ulogic;             --Dfs clocks lock signal for tiles only
signal lock_global            : std_ulogic;             --Dfs clocks lock signal for either tiles and interconnect

signal rst_ext, rst_ext_reg   : std_ulogic;             --An external reset that comes from the host computer, that triggers the system reset

--signal rst_ext_raw            : std_ulogic;             --The external reset coming out from the IO tile
--signal rst_ext_raw_sync1      : std_ulogic;             --The external reset coming out from the IO tile, first synchronizing ff
--signal rst_ext_raw_sync       : std_ulogic;             --The external reset coming out from the IO tile, second synchronizing ff
--signal counter_rst_ext        : unsigned(7 downto 0);   --A counter to automatically stop the external reset

-- NoC
signal clk_noc                : std_ulogic;--_vector(0 downto 0);        --Clock for the NoC (the output of the DFS is always a vector)
signal rstn_noc               : std_ulogic;             --Reset for the NoC
signal lock_noc               : std_ulogic;             --Lock of the NoC clock
signal noc_freq_data          : std_logic_vector(GM_FREQ_DW-1 downto 0);  --GM change: input freq data
signal noc_freq_valid         : std_logic;                                --GM change: freq data empty

-- UART
signal uart_rxd_int           : std_logic;
signal uart_txd_int           : std_logic;
signal uart_ext_addr          : std_logic_vector (CFG_UART1_FIFO-1 downto 0);
signal uart_ext_data          : std_logic_vector (CFG_UART1_FIFO-1 downto 0);
signal uart_ext_valid         : std_logic;

--signal uart_ctsn_int : std_logic;
--signal uart_rtsn_int : std_logic;
--signal uart_cts_int : std_logic;
--signal uart_rts_int : std_logic;


-- Memory bus
signal buf_ddr_ahbsi   : ahb_slv_in_vector_type(0 to CFG_NMEM_TILE-1);      --Connection between memory buffer and latency emulator
signal buf_ddr_ahbso   : ahb_slv_out_vector_type(0 to CFG_NMEM_TILE-1);

signal noc_ddr_ahbsi   : ahb_slv_in_vector_type(0 to CFG_NMEM_TILE-1);      --Connection to/from the NoC
signal noc_ddr_ahbso   : ahb_slv_out_vector_type(0 to CFG_NMEM_TILE-1);

signal mem_ddr_ahbsi   : ahb_slv_in_vector_type(0 to CFG_NMEM_TILE-1);      --Connection to/from the memory module
signal mem_ddr_ahbso   : ahb_slv_out_vector_type(0 to CFG_NMEM_TILE-1);

signal haddr_vector    : attribute_vector(0 to CFG_NMEM_TILE-1);
signal hmask_vector    : attribute_vector(0 to CFG_NMEM_TILE-1);

-- Misc
signal cpuerr        : std_ulogic;     --Error flag from the CPU


-- Avoid clock signals optimization
attribute keep : boolean;
attribute keep of clk_board : signal is true;
attribute keep of clk_sys     : signal is true;


-- MMI64  (TODO: delete these signals that are not used)
signal mon_noc          : monitor_noc_matrix(1 to 6, 0 to CFG_TILES_NUM-1);
signal mon_mem          : monitor_mem_vector(0 to CFG_NMEM_TILE + CFG_NSLM_TILE + CFG_NSLMDDR_TILE - 1);

-- Do not delete this variable - it is used by ESP's socgen python scripts
--constant CPU_FREQ : integer := 50000;

signal temp : std_logic_vector(1 downto 0);

begin

-------------------------------------------------------------------------------
-- Leds -----------------------------------------------------------------------
-------------------------------------------------------------------------------

  -- Green LED: on when bitstream is loaded
  --green_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_GREEN, '1');
  -- Red LED: on when profpga reset does not go down
  --red_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_RED, rst_board);
  -- Other LEDs: unused
  --blue_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_BLUE, '0');
  --yellow_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_YELLOW, '0');
  -- Report when program completes

  --pragma translate_off
  process(clk_board, rstn_sys)
  begin  -- process
    if rstn_sys = '1' then
      assert cpuerr = '0' report "Program Completed!" severity failure;
    end if;
  end process;
  --pragma translate_on


----------------------------------------------------------------------
--- FPGA Reset and Clock generation  ---------------------------------
----------------------------------------------------------------------

  --Board clock generation
  clk_sim: if SIMULATION = true generate
    clk_board <= clk_board_p;
  end generate clk_sim;

  clk_no_sim: if SIMULATION /= true generate
    clk_buffer_in: IBUFDS
    --generic map(
    --  CCIO_EN_M => TRUE,
    --  CCIO_EN_S => TRUE
    -- )
    port map (
      O   => clk_board,     -- 1-bit output: Buffer output
      I   => clk_board_p,   -- 1-bit input: Diff_p buffer input (connect directly to top-level port)
      IB  => clk_board_n    -- 1-bit input: Diff_n buffer input (connect directly to top-level port)
    );

  --  hbm_clk_buffer_in: IBUFDS
  --  --generic map(
  --  --  CCIO_EN_M => TRUE,
  --  --  CCIO_EN_S => TRUE
  --  -- )
  --  port map (
  --    O   => clk_hbm,     -- 1-bit output: Buffer output
  --    I   => clk_hbm_p,   -- 1-bit input: Diff_p buffer input (connect directly to top-level port)
  --    IB  => clk_hbm_n    -- 1-bit input: Diff_n buffer input (connect directly to top-level port)
  --  );
  end generate clk_no_sim;


  -- 2-stage flip-flop synchronizer for the reset
  rst_sync_in: process(clk_board)
  begin
    if rising_edge(clk_board) then
      sync_rst0 <= cpu_reset_fpga;
      sync_rst1 <= sync_rst0;
    end if;
  end process rst_sync_in;
  rst_board <= not sync_rst1;
  rstn_board <= sync_rst1;


  -- DFS for the interconnect clock
  interconnect_clock_dvfs: if CFG_HAS_DVFS /= 0 generate
    dvfs_manager_1 : clockManager
    generic map(
      PLL_FREQ => domain_freq(0),
      RANDOM_FREQ => 0
      --N_CLOCK_OUT => 1
    )
    port map(
        rst_in => rstn_init,
        clk_in => clk_sys,
        mmcm_clk_o => clk_noc,
        mmcm_locked_o => lock_noc,
        freq_data_in => noc_freq_data,
        freq_valid_in => noc_freq_valid
    );
  end generate interconnect_clock_dvfs;

  interconnect_clock_no_dvfs: if CFG_HAS_DVFS = 0 generate
    clk_noc <= clk_board;
    lock_noc <= lock_sys;
  end generate interconnect_clock_no_dvfs;

  cgi.pllctrl <= "00";
  cgi.pllrst <= rstn_board;

  --GM change: an important problem in the design of a sistem with multiple clock is that many subsystems need a synchronous reset.
  --This means that their reset must be stopped only after the locking of their clock signal, generated by the PLLs.
  --At the same time, the DFS that generates such clock signals need a reset to start its operations correctly.
  --For this reason, I decided to use two resets: the first one (the original esp reset signal for the tiles) will become the reset
  --for the local clocking resources, while my new reset (that starts after the locking of all clocks) will be the general system reset.

  --Reset for the clocking resources
  rst_clkres : rstgen         -- reset generator
  generic map (acthigh => 1, syncin => 0)
  port map (rst_board, clk_sys, lock_sys, rstn_init, open);
  lock_sys <= cgo.clklock and not rst_ext;

  --General system reset
  rst_sys : rstgen         -- reset generator
  generic map (acthigh => 1, syncin => 0)   --GM note: il segnale rst è active high, ho controllato il modulo rstgen
  port map (rst_board, clk_sys, lock_global, rstn_sys, open); --GM change: scambio rst con il mio custom
  lock_global <= lock_tiles and lock_noc and not rst_ext;

  --GM change: generate interconnect reset
  interconnect_rst: rstgen
  generic map(acthigh => 1, syncin => 0)
  port map (rst_board, clk_noc, lock_global, rstn_noc, open);


  --External reset
  --It is a reset activated by the host computer. It basically triggers the system reset, in order to restore the original state of the system.
  --It is used to reset the whole system after dynamic partial reconfiguration.

  -- The external reset runs at the frequency of clk_board. I need to convert the rst_ext_raw signal to the clk_board frequency.
  -- Note that this two-ff synchronizer works because clk_board > clk_sys.
  --external_reset_resync: process(rst_ext_raw, clk_board)
  --begin
  --if rising_edge(clk_board) then
  --  rst_ext_raw_sync1   <=   rst_ext_raw;
  --  rst_ext_raw_sync    <=   rst_ext_raw_sync1;
  --end if;
  --end process external_reset_resync;
  --
  ----Keep the external reset high for some clock cycles
  --external_reset: process(rst_board, rst_ext_raw_sync, clk_board)
  --begin
  --  if rst_board = '1' then
  --    rst_ext <= '0';
  --    counter_rst_ext <= (others => '0');
  --  elsif rising_edge(clk_board) then
  --    if rst_ext_raw_sync = '1' then
  --      rst_ext <= '1';
  --    elsif rst_ext = '1' then
  --      counter_rst_ext <= counter_rst_ext + 1;
  --      if counter_rst_ext = EXT_RST_DURATION then
  --        counter_rst_ext <= (others => '0');
  --        rst_ext <= '0';
  --      end if;
  --    end if;
  --  end if;
  --end process external_reset;

-----------------------------------------------------------------------------
-- UART pads
-----------------------------------------------------------------------------

  --uart_ctsn_int <= not uart_cts_int;
  --uart_rts_int <= not uart_rtsn_int;
  uart_rxd_pad   : inpad  generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart0_rxd, uart_rxd_int);
  uart_txd_pad   : outpad generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart0_txd, uart_txd_int);
  --uart_ctsn_pad : inpad  generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_cts, uart_cts_int);
  --uart_rtsn_pad : outpad generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_rts, uart_rts_int);

----------------------------------------------------------------------
---  DDR3 memory controller ------------------------------------------
----------------------------------------------------------------------

  --GM note: clk_sys is the 50MHz reference, compared with the clk_board which goes at 100MHz
  clkgenmigref0 : clkgen
    generic map (CFG_FABTECH, 8, 16, 0, 0, 0, 0, 0, 100000)
    port map (clk_board, clk_board, clk_sys, open, open, open, open, cgi, cgo, open, open, open);


  --gen_mig : if (SIMULATION /= true) generate

    --mig_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
    --  first_bank: if nmem = 0 generate
    --    mig_ahbram1 : ahbram
    --      generic map (
    --        hindex   => 0,
    --        tech     => 0,
    --        kbytes   => CFG_MEM_SIZE_MAIN,
    --        pipe     => 0,
    --        maccsz   => AHBDW,
    --        scantest => 0,
    --        endianness => 0
    --        )
    --      port map(
    --        rst     => rstn_noc,
    --        clk     => clk_noc,
    --        haddr   => ddr_haddr(this_ddr_index(nmem)),
    --        hmask   => ddr_hmask(this_ddr_index(nmem)),
    --        ahbsi   => mem_ddr_ahbsi(nmem),
    --        ahbso   => mem_ddr_ahbso(nmem)
    --        );
    --  end generate first_bank;
    --  generic_bank: if nmem /= 0 generate
    --    mig_ahbram1 : ahbram
    --      generic map (
    --        hindex   => 0,
    --        tech     => 0,
    --        kbytes   => CFG_MEM_SIZE_ADD,
    --        pipe     => 0,
    --        maccsz   => AHBDW,
    --        scantest => 0,
    --        endianness => 0
    --        )
    --      port map(
    --        rst     => rstn_noc,
    --        clk     => clk_noc,
    --        haddr   => ddr_haddr(this_ddr_index(nmem)),
    --        hmask   => ddr_hmask(this_ddr_index(nmem)),
    --        ahbsi   => mem_ddr_ahbsi(nmem),
    --        ahbso   => mem_ddr_ahbso(nmem)
    --        );
    --  end generate generic_bank;
    --end generate mig_loop;

   -- hbm_hconfig_gen: for nmem in 0 to CFG_NMEM_TILE-1 generate
   --   haddr_vector(nmem) <= ddr_haddr(this_ddr_index(nmem));
   --   hmask_vector(nmem) <= ddr_hmask(this_ddr_index(nmem));
   -- end generate hbm_hconfig_gen;

    hbm_i: hbm_ahb_wrapper
      generic map (
        SIMULATION  => SIMULATION,
        hindex      => 0,
        tech        => 0,
        kbytes      => 2048*1024, -- 2 GB each
        pipe        => 0,
        maccsz      => AHBDW,
        endianness  => 0,  --0 access as BE
                           --1 access as LE
        scantest    => 0
       )
      port map (
        rstn_i              => rstn_noc,
        clk_i               => clk_noc,
        hbm_clk_i           => clk_board,
        dram_stat_catrip_o  => dram_stat_catrip,
        haddr_vector_i      => ddr_haddr, --haddr_vector,
        hmask_vector_i      => ddr_hmask, --hmask_vector,
        ahbsi_i             => mem_ddr_ahbsi,
        ahbso_o             => mem_ddr_ahbso
      );
  --end generate gen_mig;

  ahbram_buffer_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
  --  --GM change: BRAM buffer instantiation
  --  ahbram_buffer_1: ahbram_buffer
  --  port map(
  --    rst_i           =>  rstn_noc,
  --    clk_i           =>  clk_noc,
  --    noc_ahbsi_i     =>  buf_ddr_ahbsi(nmem),
  --    noc_ahbso_o     =>  buf_ddr_ahbso(nmem),
  --    mem_ahbsi_o     =>  mem_ddr_ahbsi(nmem),
  --    mem_ahbso_i     =>  mem_ddr_ahbso(nmem)
  --  );
    ----GM change: latency increaser instantiation
    --ahbram_latency_simulator: ahbram_latencyIncreaser
    --generic map(
    --  LATENCY_CYCLES  =>  25
    --)
    --port map(
    --  rst_i           =>  rstn_noc,
    --  clk_i           =>  clk_noc,
    --  noc_ahbsi_i     =>  noc_ddr_ahbsi(nmem),
    --  noc_ahbso_o     =>  noc_ddr_ahbso(nmem),
    --  mem_ahbsi_o     =>  buf_ddr_ahbsi(nmem),
    --  mem_ahbso_i     =>  buf_ddr_ahbso(nmem)
    --);
    noc_ddr_ahbso(nmem) <= mem_ddr_ahbso(nmem);
    mem_ddr_ahbsi(nmem) <= noc_ddr_ahbsi(nmem);
  end generate ahbram_buffer_loop;

  --gen_mig_model : if (SIMULATION = true) generate
  --  -- pragma translate_off
  --  mig_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
  --    first_bank: if nmem = 0 generate
  --      mig_ahbram:  ahbram_sim
  --        generic map (
  --          hindex   => 0,
  --          tech     => 0,
  --          kbytes   => CFG_MEM_SIZE_MAIN,
  --          pipe     => 0,
  --          maccsz   => AHBDW,
  --          fname    => "ram.srec"
  --          )
  --        port map(
  --          rst     => rstn_noc,
  --          clk     => clk_noc,
  --          haddr   => ddr_haddr(this_ddr_index(nmem)),
  --          hmask   => ddr_hmask(this_ddr_index(nmem)),
  --          ahbsi   => mem_ddr_ahbsi(nmem),
  --          ahbso   => mem_ddr_ahbso(nmem)
  --          );
  --      end generate first_bank;
  --      generic_bank: if nmem /= 0 generate
  --        mig_ahbram:  ahbram_sim
  --        generic map (
  --          hindex   => 0,
  --          tech     => 0,
  --          kbytes   => CFG_MEM_SIZE_ADD,
  --          pipe     => 0,
  --          maccsz   => AHBDW,
  --          fname    => "ram.srec"
  --          )
  --        port map(
  --          rst     => rstn_noc,
  --          clk     => clk_noc,
  --          haddr   => ddr_haddr(this_ddr_index(nmem)),
  --          hmask   => ddr_hmask(this_ddr_index(nmem)),
  --          ahbsi   => mem_ddr_ahbsi(nmem),
  --          ahbso   => mem_ddr_ahbso(nmem)
  --          );
  --      end generate generic_bank;
  --  end generate mig_loop;
--
  --  -- pragma translate_on
  --end generate gen_mig_model;

  -----------------------------------------------------------------------------
  -- External UART
  -----------------------------------------------------------------------------
  -- I need a UART receiver external to the NoC, to manage the system reset

  external_uart: ext_uart
  generic map (
    BAUDRATE            => BAUDRATE,
    CLOCK_FREQ          => BOARD_CLOCK_FREQ,
    DATA_BYTES          => CFG_UART1_FIFO/8,
    ADDR_BYTES          => CFG_UART1_FIFO/8
  )
  port map(
    clk_i               => clk_board,
    rst_i               => rst_board,
    addr_o              => uart_ext_addr,
    data_o              => uart_ext_data,
    valid_o             => uart_ext_valid,
    rx                  => uart_rxd_int
  );

  external_reset: process (clk_board, cpu_reset_fpga)
  begin
    if cpu_reset_fpga = '0' then
        rst_ext_reg <= '0';
    elsif rising_edge(clk_board) then
      if uart_ext_valid = '1' and uart_ext_addr = x"600003FC" then
        rst_ext_reg <= uart_ext_data(0);
      end if;
    end if;
  end process;
  rst_ext <= rst_ext_reg;
  -----------------------------------------------------------------------------
  -- ESP
  -----------------------------------------------------------------------------

  esp_1: esp
    generic map (
      SIMULATION             => SIMULATION)
    port map (
      rstn_sys               => rstn_sys,
      rstn_init              => rstn_init,
      clk_sys                => clk_sys,
      clk_noc                => clk_noc,
      rstn_noc               => rstn_noc,
      pllbypass              => (others => '0'),
      lock_tiles             => lock_tiles,
      uart_rxd               => uart_rxd_int,
      uart_txd               => uart_txd_int,
      uart_ctsn              => '1',
      uart_rtsn              => open,
      cpuerr                 => cpuerr,
      ddr_ahbsi              => noc_ddr_ahbsi,
      ddr_ahbso              => noc_ddr_ahbso,
      -- Monitor signals
      mon_noc                => mon_noc,
      mon_mem                => mon_mem,
      rst_ext_out            => open,
      freq_data_out          => noc_freq_data,  --GM change: input freq data
      freq_valid_out         => noc_freq_valid --GM change: freq data empty
      );

end;


