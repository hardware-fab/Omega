-- Copyright (c) 2011-2023 Columbia University, System Level Design Group
-- SPDX-License-Identifier: Apache-2.0

------------------------------------------------------------------------------
--  ESP - profpga - TA1 - xc7v2000t
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
       
        
use work.grlib_config.all;
use work.amba.all;
use work.stdlib.all;
use work.devices.all;
use work.gencomp.all;
use work.leon3.all;
use work.uart.all;
use work.misc.all;
use work.net.all;
use work.svga_pkg.all;
library unisim;
-- pragma translate_off
use work.sim.all;
-- pragma translate_on
use unisim.VCOMPONENTS.all;
use work.monitor_pkg.all;
use work.sldacc.all;
use work.tile.all;
use work.nocpackage.all;
use work.cachepackage.all;
use work.coretypes.all;
use work.config.all;
use work.esp_global.all;
use work.socmap.all;
use work.tiles_pkg.all;

use work.esp_csr_pkg.all; --GM change: I need this library for freq data info

entity top is
  generic (
    SIMULATION          : boolean := false
  );
  port (
    clk_board_p           : in  std_ulogic;  -- 100 MHz clock
    clk_board_n           : in  std_ulogic;  -- 100 MHz clock
    profpga_sync0_p       : in  std_ulogic;
    profpga_sync0_n       : in  std_ulogic;
    reset                 : in    std_ulogic;
    uart_rxd              : in    std_ulogic;
    uart_txd              : out   std_ulogic;
    uart_cts              : in    std_ulogic;
    uart_rts              : out   std_ulogic;
    LED_RED               : out   std_ulogic;
    LED_GREEN             : out   std_ulogic;
    LED_BLUE              : out   std_ulogic;
    LED_YELLOW            : out   std_ulogic
   );
end;


architecture rtl of top is

--GM change: aggiungo il modulo che genera il reset
component profpga_clocksync is
  generic (
    CLK_CORE_COMPENSATION : string := "DELAYED" -- "DELAYED" , "DELAYED_XVUS" or "ZHOLD"
  );
  port (
    -- access to FPGA pins
    clk_p           : in  std_ulogic;
    clk_n           : in  std_ulogic;
    sync_p          : in  std_ulogic;
    sync_n          : in  std_ulogic;
    -- clock from pad
    clk_o           : out std_ulogic;
    -- clock feedback (either clk_o or 1:1 output from MMCM/PLL)
    clk_i           : in  std_ulogic;
    clk_locked_i    : in  std_ulogic;
    -- configuration access from profpga_infrastructure
    mmi64_clk       : in  std_ulogic;
    mmi64_reset     : in  std_ulogic;
    cfg_dn_i        : in  std_ulogic_vector(19 downto 0);
    cfg_up_o        : out std_ulogic_vector(19 downto 0);
    -- sync events
    user_reset_o    : out std_ulogic;
    user_strobe1_o  : out std_ulogic;
    user_strobe2_o  : out std_ulogic;
    user_event_id_o : out std_ulogic_vector(7 downto 0);
    user_event_en_o : out std_ulogic
  );
end component profpga_clocksync;
  
--GM change: I add the declaration of the DFS module
component clockManager
  generic(
    PLL_FREQ                                 :    integer := 1;
    RANDOM_FREQ                              :    integer := 0;
    N_CLOCK_OUT                              :    integer := 1
  );
  port (
    rst_in                                   :     in std_logic;
    clk_in                                   :     in std_logic;
    mmcm_clk_o                               :     out std_ulogic_vector(N_CLOCK_OUT-1 downto 0);
    mmcm_locked_o                            :     out std_logic;
    freq_data_in                             :     in std_logic_vector(8-1 downto 0);
    freq_valid_in                            :     in std_logic
    );
end component;

function set_ddr_index (
  constant n : integer range 0 to 3)
  return integer is
begin
  if n > (MEM_ID_RANGE_MSB) then
    return MEM_ID_RANGE_MSB;
  else
    return n;
  end if;
end set_ddr_index;

constant this_ddr_index : attribute_vector(0 to 3) := (
  0 => set_ddr_index(0),
  1 => set_ddr_index(1),
  2 => set_ddr_index(2),
  3 => set_ddr_index(3)
  );

--Duration of the external reset pulse
constant EXT_RST_DURATION : integer := 100;

-------------------------------------------------------------------------------
-- Signals --------------------------------------------------------------------
-------------------------------------------------------------------------------

-- Clock and reset
signal rst_sim            : std_ulogic;             --Input reset (used only in simulation)
signal clk_board          : std_ulogic;             --Clock generated by profpga_clocksync. Freq: 100MHz
signal rst_profpga        : std_ulogic;             --Reset generated by profpga_clocksync.

signal clk_sys            : std_ulogic;             --Main system clock sent to the tiles
signal lock_sys           : std_ulogic;             --Lock signal of the main system clock

signal rstn_profpga       : std_ulogic;             --Negated profpga reset, synchronized with system clock
signal rstn_sys           : std_ulogic;             --Active low main system reset
signal rstn_init          : std_ulogic;             --Active low reset for clocking resources (synchronized with system clock)

signal cgi                : clkgen_in_type;         --Clock generator input signal for the system clock
signal cgo                : clkgen_out_type;        --Clock generator output signal for the system clock

signal lock_tiles         : std_ulogic;             --Dfs clocks lock signal for tiles only
signal lock_global        : std_ulogic;             --Dfs clocks lock signal for either tiles and interconnect

signal rst_ext            : std_ulogic;             --An external reset that comes from the host computer, that triggers the system reset
signal rst_ext_raw        : std_ulogic;             --The external reset coming out from the IO tile
signal rst_ext_raw_sync1  : std_ulogic;             --The external reset coming out from the IO tile, first synchronizing ff
signal rst_ext_raw_sync   : std_ulogic;             --The external reset coming out from the IO tile, second synchronizing ff
signal counter_rst_ext    : unsigned(7 downto 0);   --A counter to automatically stop the external reset

-- NoC
signal clk_noc            : std_ulogic_vector(0 downto 0);        --Clock for the NoC (the output of the DFS is always a vector)
signal rstn_noc           : std_ulogic;             --Reset for the NoC
signal lock_noc           : std_ulogic;             --Lock of the NoC clock
signal noc_freq_data      : std_logic_vector(GM_FREQ_DW-1 downto 0);  --GM change: input freq data
signal noc_freq_valid     : std_logic;                                --GM change: freq data empty

-- UART
signal uart_rxd_int  : std_logic;
signal uart_txd_int  : std_logic;
signal uart_ctsn_int : std_logic;
signal uart_rtsn_int : std_logic;
signal uart_cts_int : std_logic;
signal uart_rts_int : std_logic;


-- Memory bus
signal buf_ddr_ahbsi   : ahb_slv_in_vector_type(0 to MEM_ID_RANGE_MSB);      --Connection between memory buffer and latency simulator
signal buf_ddr_ahbso   : ahb_slv_out_vector_type(0 to MEM_ID_RANGE_MSB);

signal noc_ddr_ahbsi   : ahb_slv_in_vector_type(0 to MEM_ID_RANGE_MSB);      --Connection to/from the NoC
signal noc_ddr_ahbso   : ahb_slv_out_vector_type(0 to MEM_ID_RANGE_MSB);

signal mem_ddr_ahbsi   : ahb_slv_in_vector_type(0 to MEM_ID_RANGE_MSB);      --Connection to/from the memory module
signal mem_ddr_ahbso   : ahb_slv_out_vector_type(0 to MEM_ID_RANGE_MSB);


-- Misc
signal cpuerr        : std_ulogic;     --Error flag from the CPU


-- Avoid clock signals optimization
attribute keep : boolean;
attribute keep of clk_board : signal is true;
attribute keep of clk_sys     : signal is true;


-- MMI64  (TODO: delete these signals that are not used)
signal mon_ddr          : monitor_ddr_vector(0 to MEM_ID_RANGE_MSB);
signal mon_noc          : monitor_noc_matrix(1 to 6, 0 to CFG_TILES_NUM-1);
signal mon_noc_actual   : monitor_noc_matrix(0 to 1, 0 to CFG_TILES_NUM-1);
signal mon_mem          : monitor_mem_vector(0 to CFG_NMEM_TILE + CFG_NSLM_TILE + CFG_NSLMDDR_TILE - 1);
signal mon_l2           : monitor_cache_vector(0 to relu(CFG_NL2 - 1));
signal mon_llc          : monitor_cache_vector(0 to relu(CFG_NLLC - 1));
signal mon_acc          : monitor_acc_vector(0 to relu(accelerators_num-1));
signal mon_dvfs         : monitor_dvfs_vector(0 to CFG_TILES_NUM-1);

--GM: Do not delete this variable - it is used by ESP's socgen python scripts
--constant CPU_FREQ : integer := 50000;

signal temp : std_logic_vector(1 downto 0);

begin

-------------------------------------------------------------------------------
-- Leds -----------------------------------------------------------------------
-------------------------------------------------------------------------------

  -- Green LED: on when bitstream is loaded
  green_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_GREEN, '1');
  -- Red LED: on when profpga reset does not go down
  red_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_RED, rst_profpga);
  -- Other LEDs: unused
  blue_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_BLUE, '0');
  yellow_led_pad : outpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (LED_YELLOW, '0');
  -- Report when program completes
  --pragma translate_off
  process(clk_board, rstn_sys)
  begin  -- process
    if rstn_sys = '1' then
      assert cpuerr = '0' report "Program Completed!" severity failure;
    end if;
  end process;
  --pragma translate_on
    

----------------------------------------------------------------------
--- FPGA Reset and Clock generation  ---------------------------------
----------------------------------------------------------------------
  interconnect_clock_dvfs: if CFG_HAS_DVFS /= 0 generate
    dvfs_manager_1 : clockManager
    generic map(
      PLL_FREQ => domain_freq(0),
      RANDOM_FREQ => 0,
      N_CLOCK_OUT => 1
    )
    port map(
        rst_in => rstn_init,
        clk_in => clk_sys,
        mmcm_clk_o => clk_noc,
        mmcm_locked_o => lock_noc,
        freq_data_in => noc_freq_data,
        freq_valid_in => noc_freq_valid
    );
  end generate interconnect_clock_dvfs;

  interconnect_clock_no_dvfs: if CFG_HAS_DVFS = 0 generate
    clk_noc(0) <= clk_board;
    lock_noc <= lock_sys;
  end generate interconnect_clock_no_dvfs;

  cgi.pllctrl <= "00";
  cgi.pllrst <= rstn_profpga;

  --GM change: an important problem in the design of a sistem with multiple clock is that many subsystems need a synchronous reset.
  --This means that their reset must be stopped only after the locking of their clock signal, generated by the PLLs.
  --At the same time, the DFS that generates such clock signals need a reset to start its operations correctly.
  --For this reason, I decided to use two resets: the first one (the original esp reset signal for the tiles) will become the reset
  --for the local clocking resources, while my new reset (that starts after the locking of all clocks) will be the general system reset.
  reset_pad : inpad generic map (tech => CFG_FABTECH, level => cmos, voltage => x18v) port map (reset, rst_sim);

  --Reset for the clocking resources
  rst_clkres : rstgen         -- reset generator
  generic map (acthigh => 1, syncin => 0)
  port map (rst_profpga, clk_sys, lock_sys, rstn_init, open);
  lock_sys <= cgo.clklock and not rst_ext;

  --General system reset
  rst_sys : rstgen         -- reset generator
  generic map (acthigh => 1, syncin => 0)   --GM note: il segnale rst è active high, ho controllato il modulo rstgen
  port map (rst_profpga, clk_sys, lock_global, rstn_sys, rstn_profpga); --GM change: scambio rst con il mio custom
  lock_global <= lock_tiles and lock_noc and not rst_ext;
  
  --GM change: generate interconnect reset
  interconnect_rst: rstgen
  generic map(acthigh => 1, syncin => 0)
  port map (rst_profpga, clk_noc(0), lock_global, rstn_noc, open);


  --External reset
  --It is a reset activated by the host computer. It basically triggers the system reset, in order to restore the original state of the system.
  --It is used to reset the whole system after dynamic partial reconfiguration.

  -- The external reset runs at the frequency of clk_sys. I need to convert the rst_ext_raw signal to the clk_board frequency.
  -- Note that this two-ff synchronizer works because clk_board > clk_sys.
  external_reset_resync: process(rst_ext_raw, clk_board)
  begin
  if rising_edge(clk_board) then
    rst_ext_raw_sync1   <=   rst_ext_raw;
    rst_ext_raw_sync    <=   rst_ext_raw_sync1;
  end if;
  end process external_reset_resync;

  --Keep the external reset high for some clock cycles
  external_reset: process(rst_profpga, rst_ext_raw_sync, clk_board)
  begin
    if rst_profpga = '1' then
      rst_ext <= '0';
      counter_rst_ext <= (others => '0');
    elsif rst_ext_raw_sync = '1' then
      rst_ext <= '1';
    elsif rising_edge(clk_sys) then
      if rst_ext = '1' then
        counter_rst_ext <= counter_rst_ext + 1;
        if counter_rst_ext = EXT_RST_DURATION then
          counter_rst_ext <= (others => '0');
          rst_ext <= '0';
        end if;
      end if;
    end if;
  end process external_reset;

-----------------------------------------------------------------------------
-- UART pads
-----------------------------------------------------------------------------

  uart_ctsn_int <= not uart_cts_int;
  uart_rts_int <= not uart_rtsn_int;
  uart_rxd_pad   : inpad  generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_rxd, uart_rxd_int);
  uart_txd_pad   : outpad generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_txd, uart_txd_int);
  uart_ctsn_pad : inpad  generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_cts, uart_cts_int);
  uart_rtsn_pad : outpad generic map (level => cmos, voltage => x18v, tech => CFG_FABTECH) port map (uart_rts, uart_rts_int);

----------------------------------------------------------------------
---  DDR3 memory controller ------------------------------------------
----------------------------------------------------------------------

  --GM note: clk_sys is the 50MHz reference, compared with the clk_board which goes at 100MHz
  clkgenmigref0 : clkgen
    generic map (CFG_FABTECH, 16, 32, 0, 0, 0, 0, 0, 100000)
    port map (clk_board, clk_board, clk_sys, open, open, open, open, cgi, cgo, open, open, open);


  gen_mig : if (SIMULATION /= true) generate

    mig_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
      first_bank: if nmem = 0 generate
        mig_ahbram1 : ahbram
          generic map (
            hindex   => 0,
            tech     => 0,
            kbytes   => CFG_MEM_SIZE_MAIN,
            pipe     => 0,
            maccsz   => AHBDW,
            scantest => 0,
            endianness => 0
            )
          port map(
            rst     => rstn_noc,
            clk     => clk_noc(0),
            haddr   => ddr_haddr(this_ddr_index(nmem)),
            hmask   => ddr_hmask(this_ddr_index(nmem)),
            ahbsi   => mem_ddr_ahbsi(nmem),
            ahbso   => mem_ddr_ahbso(nmem)
            );
      end generate first_bank;
      generic_bank: if nmem /= 0 generate
        mig_ahbram1 : ahbram
          generic map (
            hindex   => 0,
            tech     => 0,
            kbytes   => CFG_MEM_SIZE_ADD,
            pipe     => 0,
            maccsz   => AHBDW,
            scantest => 0,
            endianness => 0
            )
          port map(
            rst     => rstn_noc,
            clk     => clk_noc(0),
            haddr   => ddr_haddr(this_ddr_index(nmem)),
            hmask   => ddr_hmask(this_ddr_index(nmem)),
            ahbsi   => mem_ddr_ahbsi(nmem),
            ahbso   => mem_ddr_ahbso(nmem)
            );
      end generate generic_bank;
    end generate mig_loop;

    --GM change: genero il reset con il clock sync
    clocksync: profpga_clocksync
      port map(

      clk_p            => clk_board_p,
      clk_n            => clk_board_n,
      sync_p           => profpga_sync0_p,
      sync_n           => profpga_sync0_n,
      clk_o            => clk_board,
      clk_i            => clk_board,
      clk_locked_i     => '1',
      mmi64_clk        => '0',
      mmi64_reset      => '0',
      cfg_dn_i         => (others => '0'),
      cfg_up_o         => open,
      user_reset_o     => rst_profpga,
      user_strobe1_o   => open,
      user_strobe2_o   => open,
      user_event_id_o  => open,
      user_event_en_o  => open
      );

  end generate gen_mig;

  ahbram_buffer_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
    --GM change: BRAM buffer instantiation
    ahbram_buffer_1: ahbram_buffer
    port map(
      rst_i           =>  rstn_noc,
      clk_i           =>  clk_noc(0),
      noc_ahbsi_i     =>  buf_ddr_ahbsi(nmem),
      noc_ahbso_o     =>  buf_ddr_ahbso(nmem),
      mem_ahbsi_o     =>  mem_ddr_ahbsi(nmem),
      mem_ahbso_i     =>  mem_ddr_ahbso(nmem)
    );
    --GM change: latency increaser instantiation
    ahbram_latency_simulator: ahbram_latencyIncreaser
    generic map(
      LATENCY_CYCLES  =>  25
    )
    port map(
      rst_i           =>  rstn_noc,
      clk_i           =>  clk_noc(0),
      noc_ahbsi_i     =>  noc_ddr_ahbsi(nmem),
      noc_ahbso_o     =>  noc_ddr_ahbso(nmem),
      mem_ahbsi_o     =>  buf_ddr_ahbsi(nmem),
      mem_ahbso_i     =>  buf_ddr_ahbso(nmem)
    );
  end generate ahbram_buffer_loop;

  gen_mig_model : if (SIMULATION = true) generate
    -- pragma translate_off
    rst_profpga <= rst_sim;     --GM change: adding this for simulation. Don't know how it worked without this!

    mig_loop: for nmem in 0 to CFG_NMEM_TILE-1 generate
      first_bank: if nmem = 0 generate
        mig_ahbram:  ahbram_sim
          generic map (
            hindex   => 0,
            tech     => 0,
            kbytes   => CFG_MEM_SIZE_MAIN,
            pipe     => 0,
            maccsz   => AHBDW,
            fname    => "ram.srec"
            )
          port map(
            rst     => rstn_noc,
            clk     => clk_noc(0),
            haddr   => ddr_haddr(this_ddr_index(nmem)),
            hmask   => ddr_hmask(this_ddr_index(nmem)),
            ahbsi   => mem_ddr_ahbsi(nmem),
            ahbso   => mem_ddr_ahbso(nmem)
            );
        end generate first_bank;
        generic_bank: if nmem /= 0 generate
          mig_ahbram:  ahbram_sim
          generic map (
            hindex   => 0,
            tech     => 0,
            kbytes   => CFG_MEM_SIZE_ADD,
            pipe     => 0,
            maccsz   => AHBDW,
            fname    => "ram.srec"
            )
          port map(
            rst     => rstn_noc,
            clk     => clk_noc(0),
            haddr   => ddr_haddr(this_ddr_index(nmem)),
            hmask   => ddr_hmask(this_ddr_index(nmem)),
            ahbsi   => mem_ddr_ahbsi(nmem),
            ahbso   => mem_ddr_ahbso(nmem)
            );
        end generate generic_bank;
    end generate mig_loop;

    clk_board <= clk_board_p;

    -- pragma translate_on
  end generate gen_mig_model;

  -----------------------------------------------------------------------------
  -- ESP
  -----------------------------------------------------------------------------

  esp_1: esp
    generic map (
      SIMULATION             => SIMULATION)
    port map (
      rstn_sys               => rstn_sys,
      rstn_init              => rstn_init,
      clk_sys                => clk_sys,
      clk_noc                => clk_noc(0),
      rstn_noc               => rstn_noc,
      pllbypass              => (others => '0'),
      lock_tiles             => lock_tiles,
      uart_rxd               => uart_rxd_int,
      uart_txd               => uart_txd_int,
      uart_ctsn              => uart_ctsn_int,
      uart_rtsn              => uart_rtsn_int,
      cpuerr                 => cpuerr,
      ddr_ahbsi              => noc_ddr_ahbsi,
      ddr_ahbso              => noc_ddr_ahbso,
      -- Monitor signals
      mon_noc                => mon_noc,
      mon_acc                => mon_acc,
      mon_mem                => mon_mem,
      mon_l2                 => mon_l2,
      mon_llc                => mon_llc,
      mon_dvfs               => mon_dvfs,
      rst_ext_out            => rst_ext_raw,
      freq_data_out          => noc_freq_data,  --GM change: input freq data
      freq_valid_out         => noc_freq_valid --GM change: freq data empty
      );

end;


