------------------------------------------------------------------------------
--  This file is a part of the VESPA SoC Prototyping Framework
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the Apache 2.0 License.
--
-- File:    dual_clock_fifo_pkg.vhd
-- Authors: Gabriele Montanaro
--          Andrea Galimberti
--          Davide Zoni
-- Company: Politecnico di Milano
-- Mail:    name.surname@polimi.it
--
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package dual_clock_fifo_pkg is

--component dual_clock_fifo0
--    generic (
--      depth : integer;
--      width : integer);
--    port (
--      clk      : in  std_logic;
--      rst      : in  std_logic;
--      rdreq    : in  std_logic;
--      wrreq    : in  std_logic;
--      data_in  : in  std_logic_vector(width-1 downto 0);
--      empty    : out std_logic;
--      full     : out std_logic;
--      data_out : out std_logic_vector(width-1 downto 0));
--end component;

end dual_clock_fifo_pkg;
