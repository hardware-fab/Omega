package sim_uart_pkg;

    // UART_CLK_DIV_DEF           = clk / (16 * baud_rate)
    // SIM_UART_NUM_CLK_TICKS_BIT = clk / baud_rate


// BaudRate 1000000 bit/s @ 50MHz

    //parameter UART_CLK_DIV_DEF 				=	8'd3; 
	//parameter SIM_HALF_CLK_PERIOD_DEF       =	10; 
	//parameter SIM_UART_NUM_CLK_TICKS_BIT    =	50;

// BaudRate 115200 bit/s @ 50MHz

    //parameter UART_CLK_DIV_DEF 				=	8'd27; 
	//parameter SIM_HALF_CLK_PERIOD_DEF       =	10; 
	//parameter SIM_UART_NUM_CLK_TICKS_BIT    =	434;
	
// BaudRate 38400 bit/s @ 100MHz
   parameter UART_CLK_DIV_DEF              =   8'd163;
   parameter SIM_HALF_CLK_PERIOD_DEF       =   5;
   parameter SIM_UART_NUM_CLK_TICKS_BIT    =   2604;


// BaudRate 38400 bit/s @ 50MHz
//    parameter UART_CLK_DIV_DEF              =   8'd81;
//    parameter SIM_HALF_CLK_PERIOD_DEF       =   10;
//    parameter SIM_UART_NUM_CLK_TICKS_BIT    =   1302;



    parameter UART_NUM_CLK_TICKS_BIT 		= SIM_UART_NUM_CLK_TICKS_BIT;
    parameter UART_NUM_DWORD_BITS			= 8;
	parameter UART_NUM_STOP_BITS			= 1;
endpackage
 
