//----------------------------------------------------------------------------
//  This file is a part of the VESPA SoC Prototyping Framework
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the Apache 2.0 License.
//
// File:    bram18_old.vhd
// Authors: Gabriele Montanaro
//          Andrea Galimberti
//          Davide Zoni
// Company: Politecnico di Milano
// Mail:    name.surname@polimi.it
//
// ----------------------------------------------------------------------------

module bram18 #(
    parameter READ_WIDTH            = 18,
    parameter WRITE_WIDTH           = 18,
    parameter ADDR_WIDTH            = 10,
    parameter WE_WIDTH              = 2
    )
    (
    input                        clk,
    input                        reset,
    input  [ADDR_WIDTH-1:0]      addr_i,
    input                        valid_i,
    output [READ_WIDTH-1:0]      data_o
    );
    wire [WRITE_WIDTH-1:0] data_i ;
    wire [WE_WIDTH-1:0]    we ;
    wire                   regce;
    assign  we      = { WE_WIDTH{1'b0}    };
    assign  data_i  = { WRITE_WIDTH{1'b0} };
    assign  regce   = 1'b0;
    BRAM_SINGLE_MACRO #(
        .BRAM_SIZE("18Kb"), // Target BRAM, "18Kb" or "36Kb" 
        .DEVICE("7SERIES"), // Target Device: "7SERIES" 
        .DO_REG(0), // Optional output register (0 or 1)
        .INIT(18'b000000000000000000), // Initial values on output port
        .INIT_FILE ("NONE"),
        .WRITE_WIDTH(WRITE_WIDTH), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .READ_WIDTH(READ_WIDTH),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        .SRVAL(18'b000000000000000000), // Set/Reset value for port output
        .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
        .INIT_00(256'h1e001e001d001d001cc01c001b001b001ae01a001900190014000f000a000500),
.INIT_01(256'h23c023a023802360236023202300230022e0220021202100200020001f001f00),
.INIT_02(256'h24e024a024a02480246024402400240023e023c023a023602360234023002300),
.INIT_03(256'h250025a025a0258025402520250024e024c024c024a024802440242024202400),
.INIT_04(256'h26e026c026802680266026202620260025c025c0258025802540252025202500),
.INIT_05(256'h27c027c027a0276027402740272026e026e026a02680268026402620260026e0),
.INIT_06(256'h28c028a028802880288028002800280028002800276027602760272027202700),
.INIT_07(256'h29c029c029c02960294029402920290028e028a028a0288028402840282028e0),
.INIT_08(256'h2ac02aa02aa02a802a602a202a002a0029e029a02980296029402920292029e0),
.INIT_09(256'h2be02ba02b802b802b402b402b202b202aa02aa02aa02a602a602a402a002a00),
.INIT_0A(256'h2ce02ce02c802c802c402c202c202c002be02bc02b802b802b402b402b202be0),
.INIT_0B(256'h2de02da02da02d602d602d202d202d002cc02cc02c802c802c602c202c202ce0),
.INIT_0C(256'h2ee02ec02e802e802e402e402e002e002de02da02da02d802d602d202d002d00),
.INIT_0D(256'h2fc02fc02f802f802f402f402f002ee02ee02ec02ec02ec02e202e202e202e00),
.INIT_0E(256'h30e030e03080308030603040302030002fc02fc02f802f802f602f202f002f00),
.INIT_0F(256'h31c031c031803160316031203100310030e030a030a0308030803020302030e0),
.INIT_10(256'h32003200320032003200320032003200320032003200320031e031e031e031e0),
.INIT_11(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_12(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_13(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_14(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_15(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_16(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_17(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_18(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_19(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_1F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_20(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_21(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_22(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_23(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_24(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_25(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_26(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_27(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_28(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_29(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_2F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_30(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_31(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_32(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_33(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_34(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_35(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_36(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_37(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_38(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_39(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3A(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3B(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3C(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3D(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3E(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INIT_3F(256'h3200320032003200320032003200320032003200320032003200320032003200),
.INITP_00(256'h0000555400000555000155540000555540015555000055550000044444040400),
.INITP_01(256'h0000555400005555000155550000555500005554000055540000555500005554),
.INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)) 
        BRAM_SINGLE_MACRO_inst (
            .DO(data_o),   // Output data, width defined by READ_WIDTH parameter
            .ADDR(addr_i), // Input address, width defined by read/write port depth look at the table below
            .CLK(clk),     // 1-bit input clock
            .DI(data_i),   // Input data port, width defined by WRITE_WIDTH parameter
            .EN(valid_i),  // 1-bit input RAM enable
            .REGCE(regce), // 1-bit input output register enable
            .RST(reset),   // 1-bit input reset
            .WE(we)        // Input write enable, width defined by write port depth look at tabel below
        );
        /////////////////////////////////////////////////////////////////////
        //  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            //
        // WRITE_WIDTH |           | WRITE Depth |            |  WE Width  //
        // ============|===========|=============|============|============//
        //    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   //
        //    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   //
        //    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   //
        //    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   //
        //    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   //
        //     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   //
        //     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   //
        //     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   //
        //     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   //
        //       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   //
        //       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   //
        //       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   //
        //       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   //
        /////////////////////////////////////////////////////////////////////
        
 endmodule
